package contants is

    constant DB_WIDTH: integer := 16;

end package contants ;