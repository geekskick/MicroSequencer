package alu_commands is
        type alu_commands_t is (alu_add1, alu_sub1, alu_inac1, alu_clac1, alu_and1, alu_or1, alu_not1, alu_xor1, alu_op2_thru, alu_lshift, alu_rshift, alu_dont_care);
end package alu_commands;
