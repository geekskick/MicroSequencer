package constants is

    constant DB_WIDTH: integer := 16;
	constant ALU_CMD_WIDTH : integer := 4;

end package constants;