-- Code your testbench here
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
port( addr: in std_logic_vector(5 downto 0);
	output: out std_logic_vector(20 downto 0)
);
end entity;

architecture struct of rom is

    -- conditions 
    -- 1  11
    -- Z  00  
    -- nZ 01
    -- xx 10

    -- branch types
    -- JUMP 00
    -- MAP  10  
    -- CALL 01
    -- RET  11


	--  M1           M2        M3      ALU 
-- NOP   000    NOP   000   NOP 0   NOP     0000
-- ARIN  001	 PCIN  001   DRM 1	PLUS    0001					
-- ARDT  010    PCDT  010
-- ARPC  011    IRDR  011           MINU    0010
-- TRDR  100    RAC	 100
-- ERROR 101    MDR   101           ACIN    0011
-- ACR   110    DRAC  110           ACZO    0100
-- ACDR  111    ZALU  111           AND     0101
--                                  OR      0110
--                                  NOT     0111
--                                  XOR     1000
--                                  THRU    1001
--                                  THRU    1010
--                                  LSHIFT  1011
--                                  RSHIFT  1100                          

type mem is array (0 to 63) of std_logic_vector(20 downto 0); 
constant microcode : mem := ( 
--location => bt & condition & M1 & M2 & M3 & next address
0 => "00" & "11" & "000" & "000" & "0" & "0000" & "000001",     -- NOP
1 => "00" & "11" & "011" & "000" & "0" & "0000" & "000111",     -- FETCH1
2 => "01" & "11" & "000" & "000" & "0" & "0000" & "010011",     -- LDAC0
3 => "00" & "11" & "000" & "000" & "1" & "0000" & "011001",     -- LDAC4
4 => "01" & "11" & "000" & "000" & "0" & "0000" & "010011",     -- STAC0
5 => "00" & "11" & "000" & "110" & "0" & "0000" & "011011",     -- STAC4
6 => "00" & "11" & "000" & "100" & "0" & "0000" & "000001",     -- MVAC1
7 => "00" & "11" & "000" & "001" & "1" & "0000" & "001001",     -- FETCH2
8 => "00" & "11" & "110" & "111" & "0" & "1001" & "000001",     -- MOVR1
9 => "10" & "10" & "011" & "011" & "0" & "0000" & "011111",     -- FETCH3
10 => "00" & "11" & "001" & "000" & "1" & "0000" & "001011",     -- JUMP1
11 => "00" & "11" & "100" & "000" & "1" & "0000" & "010001",     -- JUMP2
12 => "00" & "00" & "000" & "000" & "0" & "0000" & "001010",     -- JMPZ1
13 => "00" & "11" & "000" & "001" & "0" & "0000" & "011101",     -- NJMP1
14 => "00" & "01" & "000" & "000" & "0" & "0000" & "001010",     -- JMPNZ1
15 => "00" & "11" & "000" & "001" & "0" & "0000" & "011101",     -- JMPNZN1
16 => "00" & "11" & "000" & "111" & "0" & "0001" & "000001",     -- ADD1
17 => "00" & "11" & "000" & "010" & "0" & "0000" & "000001",     -- JUMP3
18 => "00" & "11" & "000" & "111" & "0" & "0010" & "000001",     -- SUB1
19 => "00" & "11" & "001" & "001" & "1" & "0000" & "010101",     -- STLD1
20 => "00" & "11" & "000" & "111" & "0" & "0011" & "000001",     -- INAC1
21 => "00" & "11" & "100" & "001" & "1" & "0000" & "010111",     -- STLD2
22 => "00" & "11" & "000" & "111" & "0" & "0100" & "000001",     -- CLAC1
23 => "11" & "10" & "010" & "000" & "0" & "0000" & "011111",     -- STLD3
24 => "00" & "11" & "000" & "111" & "0" & "0101" & "000001",     -- AND1
25 => "00" & "11" & "111" & "111" & "0" & "1001" & "000001",     -- LDAC5
26 => "00" & "11" & "000" & "111" & "0" & "0110" & "000001",     -- OR1
27 => "00" & "11" & "000" & "101" & "0" & "0000" & "000001",     -- STAC5
28 => "00" & "11" & "000" & "111" & "0" & "1000" & "000001",     -- XOR1
29 => "00" & "11" & "000" & "001" & "0" & "0000" & "000001",     -- NJMP2
30 => "00" & "11" & "000" & "111" & "0" & "0111" & "000001",     -- NOT1
31 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
32 => "00" & "11" & "000" & "111" & "0" & "1011" & "000001",     -- LSHIFT
33 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
34 => "00" & "11" & "000" & "111" & "0" & "1100" & "000001",     -- RSHIFT
35 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
36 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
37 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
38 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
39 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
40 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
41 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
42 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
43 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
44 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
45 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
46 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
47 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
48 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
49 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
50 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
51 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
52 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
53 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
54 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
55 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
56 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
57 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
58 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
59 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
60 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
61 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
62 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111",     -- ERROR
63 => "00" & "11" & "101" & "000" & "0" & "0000" & "011111"      -- ERROR
);  


begin

output <= microcode(to_integer(unsigned(addr)));


end architecture;