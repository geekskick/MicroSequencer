package contsants is

    constant DB_WIDTH: integer := 16;

end package contsants ;