package constants is

    constant DB_WIDTH: integer := 16;

end package constants;