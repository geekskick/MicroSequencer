package cpu_constants is
    
    constant DB_WIDTH      : integer := 16;
    constant ALU_CMD_WIDTH : integer := 4;
    constant IR_WIDTH      : integer := 5;
    
end package cpu_constants;
